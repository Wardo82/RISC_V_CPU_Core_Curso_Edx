entity main_core is
  port (
    i_clock : in std_logic;
    i_reset : in std_logic;
  ) ;
end main_core;

architecture structural* of main_core is

    signal 

begin

    -- Connect everything together


end structural* ; -- structural*