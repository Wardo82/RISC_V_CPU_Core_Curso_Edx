entity turpial_core is
  port (
    i_clock : in std_logic;
    i_reset : in std_logic;
  ) ;
end turpial_core;

architecture structural* of turpial_core is

    signal 

begin

    -- Connect everything together


end structural* ; -- structural*