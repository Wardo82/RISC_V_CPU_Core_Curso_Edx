entity data_memory is
  port (    
    clock
  ) ;
end data_memory;    

architecture behavioral of data_memory is

    signal 

begin

end behavioral ; -- behavioral