entity alu is
    port(
        i_operator1 : in std_logic_vector();
        i_operator2 : in std_logic_vector();
        o_result    : out std_logic_vector();
        o_address   : out std_logic_vector();
    );
end alu;

architecture behavioral of alu is

    signal 

begin

end behavioral ; -- behavioral